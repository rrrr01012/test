module HelloVerilog;

initial 
    begin
        $display("Hello, iverilog");
        $finish;
    end

endmodule // End of HelloVerilog